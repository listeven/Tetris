`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   16:59:14 10/15/2015
// Design Name:   Verilog
// Module Name:   X:/311Lab/BitAdder/TestModule.v
// Project Name:  BitAdder
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Verilog
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TestModule;
/*
	// Inputs
	reg a;
	reg b;
	reg Cin;
	// Outputs
	wire S;
	wire C;
	/*wire C0;
	wire C1;
	wire C2;
	wire C3;*/
	/*wire B0;
	wire B1;
	wire B2;
	wire B3;
*/



/*
	// Instantiate the Unit Under Test (UUT)
	WholeAdder uut (
		.S(S),
		.C(C),
		.a(a), 
		.b(b),
		.Cin(Cin),
	);

	initial begin
		// Initialize Inputs
		a = 1;
		b = 1;
		Cin = 0;
		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      */
endmodule

